library verilog;
use verilog.vl_types.all;
entity Semaforos_Demo is
    port(
        SW              : in     vl_logic_vector(3 downto 0);
        LEDR            : out    vl_logic_vector(17 downto 0);
        LEDG            : out    vl_logic_vector(7 downto 0);
        CLOCK_50        : in     vl_logic
    );
end Semaforos_Demo;
