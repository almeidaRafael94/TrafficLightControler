library verilog;
use verilog.vl_types.all;
entity BinUDCntEnRst4_vlg_vec_tst is
end BinUDCntEnRst4_vlg_vec_tst;
