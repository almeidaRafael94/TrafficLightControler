library verilog;
use verilog.vl_types.all;
entity CounterUp_vlg_vec_tst is
end CounterUp_vlg_vec_tst;
