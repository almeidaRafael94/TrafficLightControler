library verilog;
use verilog.vl_types.all;
entity Semaforos_Demo_vlg_vec_tst is
end Semaforos_Demo_vlg_vec_tst;
